entity KS_ADDER is 
port(
	I0,I1 : in bit_vector(0 to 15);
	A     : out bit_vector(0 to 15)
	);
entity Testbench is 
end entity Testbench;

architecture tb of Testbench is 
component ALU is 
port (
	D0, D1 : in bit_vector(15 downto 0); --inputs
	
	S0, S1 : in bit; --control inputs
	A      : out bit_vector(15 downto 0); --output vector
	C,Z    : out bit; --carry bit and zero bit
	Carryo: out bit_vector(16 downto 0)
);
end component;

signal P,Q : bit_vector(15 downto 0); --inputs
signal R   : bit_vector(15 downto 0); --output
signal T1,T2 : bit; --control inputs
signal carry,zero_bit : bit; --carry out and zero bit
signal Carrytest:	 bit_vector(16 downto 0);

begin
dut_instance : ALU
port map (D0 => P, D1 => Q, S0 => T1, S1 => T2,A => R, C => carry, Z => zero_bit, Carryo=>Carrytest );

process
begin
T1 <= '0';
T2 <= '0';
P<="0010001011111010";
Q<="0010001011111010";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="0010001011111010";
Q<="0010001011111010";

wait for 5 ns;

T1 <= '1';
T2 <= '0';
P<="0010001011111010";
Q<="0010001011111010";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="0010001011111010";
Q<="0010001011111010";

wait for 5 ns;

T1 <= '0';
T2 <= '0';
P<="0111000100000111";
Q<="0101111101011101";

wait for 5 ns;


T1 <= '0';
T2 <= '1';
P<="0111000100000111";
Q<="0101111101011101";

wait for 5 ns;


T1 <= '1';
T2 <= '0';
P<="0111000100000111";
Q<="0101111101011101";

wait for 5 ns;


T1 <= '1';
T2 <= '1';
P<="0111000100000111";
Q<="0101111101011101";

wait for 5 ns;


T1 <= '0';
T2 <= '0';
P<="0110001000001111";
Q<="1111010011111100";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="0110001000001111";
Q<="1111010011111100";

wait for 5 ns;

T1 <= '1';
T2 <= '0';
P<="0110001000001111";
Q<="1111010011111100";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="0110001000001111";
Q<="1111010011111100";

wait for 5 ns;

T1 <= '0';
T2 <= '0';
P<="0000011010010111";
Q<="1110000100101010";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="0000011010010111";
Q<="1110000100101010";

wait for 5 ns;

T1 <= '1';
T2 <= '0';
P<="0000011010010111";
Q<="1110000100101010";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="0000011010010111";
Q<="1110000100101010";

wait for 5 ns;

T1 <= '0';
T2 <= '0';
P<="1010000101111011";
Q<="0010001000110101";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="1010000101111011";
Q<="0010001000110101";

wait for 5 ns;

T1 <= '1';
T2 <= '0';
P<="1010000101111011";
Q<="0010001000110101";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="1010000101111011";
Q<="0010001000110101";

wait for 5 ns;

T1 <= '0';
T2 <= '0';
P<="1101000111111010";
Q<="0101111011101000";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="1101000111111010";
Q<="0101111011101000";

wait for 5 ns;

T1 <= '1';
T2 <= '0';
P<="1101000111111010";
Q<="0101111011101000";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="1101000111111010";
Q<="0101111011101000";

wait for 5 ns;

T1 <= '0';
T2 <= '0';
P<="1100000011100000";
Q<="1101010011111101";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="1100000011100000";
Q<="1101010011111101";

wait for 5 ns;

T1 <= '1';
T2 <= '0';
P<="1100000011100000";
Q<="1101010011111101";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="1100000011100000";
Q<="1101010011111101";

wait for 5 ns;

T1 <= '0';
T2 <= '0';
P<="1000111110010001";
Q<="1000101000100111";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="1000111110010001";
Q<="1000101000100111";

wait for 5 ns;

T1 <= '1';
T2 <= '0';
P<="1000111110010001";
Q<="1000101000100111";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="1000111110010001";
Q<="1000101000100111";

wait for 5 ns;

T1 <= '0';
T2 <= '0';
P<="0000000000000000";
Q<="0000000000000000";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="0000000000000000";
Q<="0000000000000000";

wait for 5 ns;

T1 <= '1';
T2 <= '0';
P<="0000000000000000";
Q<="0000000000000000";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="0000000000000000";
Q<="0000000000000000";

wait for 5 ns;


T1 <= '0';
T2 <= '0';
P<="0000000000000000";
Q<="1111111111111111";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="0000000000000000";
Q<="1111111111111111";

wait for 5 ns;

T1 <= '1';
T2 <= '0';
P<="0000000000000000";
Q<="1111111111111111";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="0000000000000000";
Q<="1111111111111111";

wait for 5 ns;

T1 <= '0';
T2 <= '0';
P<="1111111111111111";
Q<="0000000000000000";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="1111111111111111";
Q<="0000000000000000";

wait for 5 ns;
T1 <= '1';
T2 <= '0';
P<="1111111111111111";
Q<="0000000000000000";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="1111111111111111";
Q<="0000000000000000";

wait for 5 ns;

T1 <= '0';
T2 <= '0';
P<="1111111111111111";
Q<="1111111111111111";

wait for 5 ns;

T1 <= '0';
T2 <= '1';
P<="1111111111111111";
Q<="1111111111111111";

wait for 5 ns;

T1 <= '1';
T2 <= '0';
P<="1111111111111111";
Q<="1111111111111111";

wait for 5 ns;

T1 <= '1';
T2 <= '1';
P<="1111111111111111";
Q<="1111111111111111";

wait for 5 ns;

end process;
end tb;
entity OR2 is 
port (
	E,F : in bit;
	G   : out bit	
);
end entity OR2;


architecture struct of OR2 is 
begin

G <= E OR F;

end struct ;